FROM spiceai/spiceai:latest-models
ADD spicepod.yaml /app
